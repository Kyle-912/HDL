library ieee;
use ieee.std_logic_1164.all;

entity datapath is
  generic (
    width : positive := 16);
  port (
    clk       : in  std_logic;
    rst       : in  std_logic;
    en        : in  std_logic;
    valid_in  : in  std_logic;
    valid_out : out std_logic;
    in1       : in  std_logic_vector(width - 1 downto 0);
    in2       : in  std_logic_vector(width - 1 downto 0);
    in3       : in  std_logic_vector(width - 1 downto 0);
    in4       : in  std_logic_vector(width - 1 downto 0);
    output    : out std_logic_vector(width * 2 downto 0));
end datapath;

-- TODO: Implement the structural description of the datapath shown in
-- datapath.pdf by instantiating your add_pipe and mult_pipe entities. You may
-- also use the provided reg entity, or you can create your own.

architecture STR of datapath is

begin

end STR;
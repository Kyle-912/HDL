library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use ieee.math_real.all;

entity fib_tb is
end fib_tb;

architecture tb of fib_tb is
begin

end tb;